
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DEM_00_99_HT_7DOAN is
	Port ( CKHT : in  STD_LOGIC;
			  BTN_N : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
           SSEG : out  STD_LOGIC_VECTOR (7 downto 0);
           BELL : out  STD_LOGIC;
           ANODE : OUT  STD_LOGIC_VECTOR (7 downto 0));
end DEM_00_99_HT_7DOAN;

architecture Behavioral of DEM_00_99_HT_7DOAN is
SIGNAL ENA5HZ,ENA2HZ, ENA1KHZ, RST : STD_LOGIC;
SIGNAL DONVIA,CHUCA,DONVIB,CHUCB,DONVIC,CHUCC: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL DAU_CHAM_8LED: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ENA_GIAIMA_8LED: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL BT1,BT2,BT3: STD_LOGIC;
begin
	BELL <= '1';
	RST <= NOT BTN_N(0);
	DAU_CHAM_8LED <= X"FF";
	ENA_GIAIMA_8LED <= X"DB"; 
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
			PORT MAP(	CKHT => CKHT,
							ENA5HZ => ENA5HZ,
							ENA2HZ => ENA2HZ,
							ENA1KHZ => ENA1KHZ);
DEM_1BIT_BTNA: ENTITY WORK.DEM_1BIT_BTN
		PORT MAP(	CKHT => CKHT,
						RST => RST,
						BTN => NOT BTN_N(1),
						Q => BT1);
DEM_1BIT_BTNB: ENTITY WORK.DEM_1BIT_BTN
		PORT MAP(	CKHT => CKHT,
						RST => RST,
						BTN => NOT BTN_N(2),
						Q => BT2);
DEM_1BIT_BTNC: ENTITY WORK.DEM_1BIT_BTN
		PORT MAP(	CKHT => CKHT,
						RST => RST,
						BTN => NOT BTN_N(3),
						Q => BT3);
DEM_2SOA:	ENTITY WORK.DEM_2SOA
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_DB => ENA5HZ,
							ENA_SS => BT1,
							ENA_SS1 => BT3,
							DONVI => DONVIA,
							CHUC => CHUCA); -- THEM CHO NAY
DEM_2SOB:	ENTITY WORK.DEM_2SOB
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_DB => ENA5HZ,
							ENA_SS => BT2,
							ENA_SS1 => BT3,
							DONVI => DONVIB,
							CHUC => CHUCB);							
DEM_2SOC:	ENTITY WORK.DEM_2SOC
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_DB => ENA2HZ,
							ENA_SS => BT3,
							DONVIA => DONVIA,
							CHUCA  => CHUCA,
							DONVIB => DONVIB,
							CHUCB  => CHUCB,
							DONVI => DONVIC,
							CHUC => CHUCC);


HIENTHI_2LED: ENTITY WORK.GIAIMA_HIENTHI_8LED_7DOAN
			PORT MAP(
					CKHT => CKHT,
					ENA1KHZ => ENA1KHZ,
					LED70 => DONVIA,
					LED71 => CHUCA, --- NHO SUA CHO NAY
					LED72 => X"F",
					LED73 => DONVIB,
					LED74 => CHUCB,
					LED75 => X"F",
					LED76 => DONVIC,
					LED77 => CHUCC,
					DAU_CHAM_8LED => DAU_CHAM_8LED,
					ENA_GIAIMA_8LED => ENA_GIAIMA_8LED,
					ANODE => ANODE,
					SSEG => SSEG);
end Behavioral;

