
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;


entity LCD_GAN_DULIEU_1SO_TO is
    Port ( ENA :in std_logic;
			  CH_GIO,DV_GIO,CH_PHUT,DV_PHUT,CH_GIAY,DV_GIAY,CH_ND,DV_ND : in  STD_LOGIC_VECTOR (3 downto 0);
			  LCD_CH_GIO,LCD_DV_GIO,LCD_CH_PHUT,LCD_DV_PHUT,LCD_CH_GIAY,LCD_DV_GIAY,LCD_CH_ND,LCD_DV_ND,LCD_CHU_TO : in  STD_LOGIC_VECTOR (47 downto 0);
           LCD_HANG_1 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_HANG_2 : out  STD_LOGIC_VECTOR (159 downto 0);
			  LCD_HANG_3 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_HANG_4 : out  STD_LOGIC_VECTOR (159 downto 0));
end LCD_GAN_DULIEU_1SO_TO;

architecture Behavioral of LCD_GAN_DULIEU_1SO_TO is

begin
	LCD_HANG_1( 7 DOWNTO 0) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_GIO(47 DOWNTO 40);  
	LCD_HANG_1( 15 DOWNTO 8) 	<= X"3"&CH_GIO WHEN ENA = '0' ELSE LCD_CH_GIO(39 DOWNTO 32);   
	LCD_HANG_1( 23 DOWNTO 16) 	<= X"3"&DV_GIO WHEN ENA = '0' ELSE LCD_CH_GIO(31 DOWNTO 24);  
	LCD_HANG_1( 31 DOWNTO 24) 	<= X"20" WHEN ENA = '0' ELSE LCD_DV_GIO(47 DOWNTO 40);
	LCD_HANG_1( 39 DOWNTO 32) 	<= X"20" WHEN ENA = '0' ELSE LCD_DV_GIO(39 DOWNTO 32);  
	LCD_HANG_1( 47 DOWNTO 40) 	<= X"20" WHEN ENA = '0' ELSE LCD_DV_GIO(31 DOWNTO 24);  
	LCD_HANG_1( 55 DOWNTO 48) 	<= X"20";  ---- 6 -----
	LCD_HANG_1( 63 DOWNTO 56) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_PHUT(47 DOWNTO 40); 
	LCD_HANG_1( 71 DOWNTO 64) 	<= X"3"&CH_PHUT WHEN ENA = '0' ELSE LCD_CH_PHUT(39 DOWNTO 32); 
	LCD_HANG_1( 79 DOWNTO 72) 	<= X"3"&DV_PHUT WHEN ENA = '0' ELSE LCD_CH_PHUT(31 DOWNTO 24); 
	LCD_HANG_1( 87 DOWNTO 80) 	<= X"20" WHEN ENA = '0' ELSE LCD_DV_PHUT(47 DOWNTO 40); 
	LCD_HANG_1( 95 DOWNTO 88) 	<= X"20" WHEN ENA = '0' ELSE LCD_DV_PHUT(39 DOWNTO 32);
	LCD_HANG_1( 103 DOWNTO 96)	<= X"20" WHEN ENA = '0' ELSE LCD_DV_PHUT(31 DOWNTO 24);
	LCD_HANG_1( 111 DOWNTO 104) <= X"20";
	LCD_HANG_1( 119 DOWNTO 112) <= X"20" WHEN ENA = '0' ELSE LCD_CH_GIAY(47 DOWNTO 40); 
	LCD_HANG_1( 127 DOWNTO 120) <= X"3"&CH_GIAY WHEN ENA = '0' ELSE LCD_CH_GIAY(39 DOWNTO 32); 
	LCD_HANG_1( 135 DOWNTO 128) <= X"3"&DV_GIAY WHEN ENA = '0' ELSE LCD_CH_GIAY(31 DOWNTO 24); 
	LCD_HANG_1( 143 DOWNTO 136) <= X"20" WHEN ENA = '0' ELSE LCD_DV_GIAY(47 DOWNTO 40);
	LCD_HANG_1( 151 DOWNTO 144) <= X"20" WHEN ENA = '0' ELSE LCD_DV_GIAY(39 DOWNTO 32); 
	LCD_HANG_1( 159 DOWNTO 152) <= X"20" WHEN ENA = '0' ELSE LCD_DV_GIAY(31 DOWNTO 24); 		

	LCD_HANG_2( 7 DOWNTO 0) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_GIO(23 DOWNTO 16);  
	LCD_HANG_2( 15 DOWNTO 8) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_GIO(15 DOWNTO 8); 
	LCD_HANG_2( 23 DOWNTO 16) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_GIO(7 DOWNTO 0); 
	LCD_HANG_2( 31 DOWNTO 24) 	<= X"20" WHEN ENA = '0' ELSE LCD_DV_GIO(23 DOWNTO 16); 
	LCD_HANG_2( 39 DOWNTO 32) 	<= X"20" WHEN ENA = '0' ELSE LCD_DV_GIO(15 DOWNTO 8); 
	LCD_HANG_2( 47 DOWNTO 40) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_GIO(7 DOWNTO 0); 
	LCD_HANG_2( 55 DOWNTO 48) 	<= X"20";
	LCD_HANG_2( 63 DOWNTO 56) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_PHUT(23 DOWNTO 16);  
	LCD_HANG_2( 71 DOWNTO 64) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_PHUT(15 DOWNTO 8);  
	LCD_HANG_2( 79 DOWNTO 72) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_PHUT(7 DOWNTO 0); 
	LCD_HANG_2( 87 DOWNTO 80) 	<= X"20" WHEN ENA = '0' ELSE LCD_DV_PHUT(23 DOWNTO 16); 
	LCD_HANG_2( 95 DOWNTO 88) 	<= X"20" WHEN ENA = '0' ELSE LCD_DV_PHUT(15 DOWNTO 8);
	LCD_HANG_2( 103 DOWNTO 96)	<= X"20" WHEN ENA = '0' ELSE LCD_DV_PHUT(7 DOWNTO 0);
	LCD_HANG_2( 111 DOWNTO 104) <= X"20";
	LCD_HANG_2( 119 DOWNTO 112) <= X"20" WHEN ENA = '0' ELSE LCD_CH_GIAY(23 DOWNTO 16);
	LCD_HANG_2( 127 DOWNTO 120) <= X"20" WHEN ENA = '0' ELSE LCD_CH_GIAY(15 DOWNTO 8);
	LCD_HANG_2( 135 DOWNTO 128) <= X"20" WHEN ENA = '0' ELSE LCD_CH_GIAY(7 DOWNTO 0);
	LCD_HANG_2( 143 DOWNTO 136) <= X"20" WHEN ENA = '0' ELSE LCD_DV_GIAY(23 DOWNTO 16);
	LCD_HANG_2( 151 DOWNTO 144) <= X"20" WHEN ENA = '0' ELSE LCD_DV_GIAY(15 DOWNTO 8);
	LCD_HANG_2( 159 DOWNTO 152) <= X"20" WHEN ENA = '0' ELSE LCD_DV_GIAY(7 DOWNTO 0);

	LCD_HANG_3( 7 DOWNTO 0) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS('N'),8);  ---- 0 -----
	LCD_HANG_3( 15 DOWNTO 8) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS('H'),8);  ---- 1 -----
	LCD_HANG_3( 23 DOWNTO 16) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS('I'),8);  ---- 2 -----
	LCD_HANG_3( 31 DOWNTO 24) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS('E'),8);  ---- 3 -----
	LCD_HANG_3( 39 DOWNTO 32) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS('T'),8);  ---- 4 -----
	LCD_HANG_3( 47 DOWNTO 40) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS(' '),8);  ---- 5 -----
	LCD_HANG_3( 55 DOWNTO 48) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS('D'),8);  ---- 6 -----
	LCD_HANG_3( 63 DOWNTO 56) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS('O'),8);  ---- 7 -----
	LCD_HANG_3( 71 DOWNTO 64) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS(':'),8);  ---- 8 -----
	LCD_HANG_3( 79 DOWNTO 72) 	<= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS(' '),8);  ---- 9 -----
	LCD_HANG_3( 87 DOWNTO 80) 	<= X"3"&CH_ND WHEN ENA = '0' ELSE LCD_CH_ND(47 DOWNTO 40);
	LCD_HANG_3( 95 DOWNTO 88) 	<= X"3"&DV_ND WHEN ENA = '0' ELSE LCD_CH_ND(39 DOWNTO 32);
	LCD_HANG_3( 103 DOWNTO 96)	<= X"00" WHEN ENA = '0' ELSE LCD_CH_ND(31 DOWNTO 24);
	LCD_HANG_3( 111 DOWNTO 104) <= CONV_STD_LOGIC_VECTOR  (CHARACTER'POS('C'),8) WHEN ENA = '0' ELSE LCD_DV_ND(47 DOWNTO 40);
	LCD_HANG_3( 119 DOWNTO 112) <= X"20" WHEN ENA = '0' ELSE LCD_DV_ND(39 DOWNTO 32);
	LCD_HANG_3( 127 DOWNTO 120) <= X"20" WHEN ENA = '0' ELSE LCD_DV_ND(31 DOWNTO 24);
	LCD_HANG_3( 135 DOWNTO 128) <= X"20" WHEN ENA = '0' ELSE CONV_STD_LOGIC_VECTOR  (CHARACTER'POS('O'),8);
	LCD_HANG_3( 143 DOWNTO 136) <= X"20" WHEN ENA = '0' ELSE LCD_CHU_TO(47 DOWNTO 40);
	LCD_HANG_3( 151 DOWNTO 144) <= X"20" WHEN ENA = '0' ELSE LCD_CHU_TO(39 DOWNTO 32);
	LCD_HANG_3( 159 DOWNTO 152) <= X"20" WHEN ENA = '0' ELSE LCD_CHU_TO(31 DOWNTO 24);

	LCD_HANG_4(7 DOWNTO 0) 		<= X"20";
	LCD_HANG_4(15 DOWNTO 8) 	<= X"20";
	LCD_HANG_4(23 DOWNTO 16) 	<= X"20";
	LCD_HANG_4(31 DOWNTO 24) 	<= X"20";
	LCD_HANG_4(39 DOWNTO 32) 	<= X"20";
	LCD_HANG_4(47 DOWNTO 40) 	<= X"20";
	LCD_HANG_4(55 DOWNTO 48) 	<= X"20";
	LCD_HANG_4(63 DOWNTO 56) 	<= X"20";
	LCD_HANG_4(71 DOWNTO 64) 	<= X"20";
	LCD_HANG_4(79 DOWNTO 72) 	<= X"20";
	LCD_HANG_4(87 DOWNTO 80) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_ND(23 DOWNTO 16);
	LCD_HANG_4(95 DOWNTO 88) 	<= X"20" WHEN ENA = '0' ELSE LCD_CH_ND(15 DOWNTO 8);
	LCD_HANG_4(103 DOWNTO 96)	<= X"20" WHEN ENA = '0' ELSE LCD_CH_ND(7 DOWNTO 0);
	LCD_HANG_4(111 DOWNTO 104) <= X"20" WHEN ENA = '0' ELSE LCD_DV_ND(23 DOWNTO 16);
	LCD_HANG_4(119 DOWNTO 112) <= X"20" WHEN ENA = '0' ELSE LCD_DV_ND(15 DOWNTO 8);
	LCD_HANG_4(127 DOWNTO 120) <= X"20" WHEN ENA = '0' ELSE LCD_DV_ND(7 DOWNTO 0);
	LCD_HANG_4(135 DOWNTO 128) <= X"20";
	LCD_HANG_4(143 DOWNTO 136) <= X"20" WHEN ENA = '0' ELSE LCD_CHU_TO(23 DOWNTO 16);
	LCD_HANG_4(151 DOWNTO 144) <= X"20" WHEN ENA = '0' ELSE LCD_CHU_TO(15 DOWNTO 8);
	LCD_HANG_4(159 DOWNTO 152) <= X"20" WHEN ENA = '0' ELSE LCD_CHU_TO(7 DOWNTO 0);
end Behavioral;

