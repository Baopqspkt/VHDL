----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:24:18 11/24/2018 
-- Design Name: 
-- Module Name:    LCD_GAN_DULIEU_HIENTHI - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity LCD_GAN_DULIEU_HIENTHI is
    Port ( DONVI:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  CHUC:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  ENA_DB,CHOPHEP,RST:IN STD_LOGIC;
			  LCD_HANG_1 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_HANG_2 : out  STD_LOGIC_VECTOR (159 downto 0);
			  LCD_HANG_3 : out  STD_LOGIC_VECTOR (159 downto 0);
			  LCD_HANG_4 : out  STD_LOGIC_VECTOR (159 downto 0));
end LCD_GAN_DULIEU_HIENTHI;

architecture Behavioral of LCD_GAN_DULIEU_HIENTHI is
TYPE MANG_DICH_TSP IS ARRAY(INTEGER RANGE 0 TO 39) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL HOVATEN_TSP : MANG_DICH_TSP:= ( 0 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--19
													1 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--19
													2 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--19
													3 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--19
													4 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('G'),8),--19
													5 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('U'),8),--19
													6 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('Y'),8),--19
													7 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8),--16
													8 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--16
													9 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
													10 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('V'),8),--16
													11 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8),--16
													12 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--16
													13 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
													14 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('V'),8),--16
													15 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('Y'),8),--16
													16 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
													17 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--1
													18 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--2                              
													19 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--3 
													
													20 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--4
													21 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--5
													22 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--6
													23 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--7
													24 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--8                  
													25 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--9	                                 
													26 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--10
													27 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--11
													28 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--12
													29 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--13
													30 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--14                             
													31 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--15 
													32 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--7
													33 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--8                  
													34 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--9	                                 
													35 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--10
													36 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--11
													37 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--12
													38 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--13
													39 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8)--14                              
													);
													
TYPE MANG_DICH_PST IS ARRAY(INTEGER RANGE 0 TO 39) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL HOVATEN_PST : MANG_DICH_PST:= ( 0 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--19
													1 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--19
													2 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--19
													3 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--19
													4 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('G'),8),--19
													5 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('U'),8),--19
													6 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('Y'),8),--19
													7 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8),--16
													8 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--16
													9 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
													10 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('V'),8),--16
													11 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8),--16
													12 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--16
													13 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
													14 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('V'),8),--16
													15 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('Y'),8),--16
													16 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
													17 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--1
													18 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--2                              
													19 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--3 
													
													20 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--4
													21 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--5
													22 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--6
													23 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--7
													24 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--8                  
													25 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--9	                                 
													26 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--10
													27 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--11
													28 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--12
													29 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--13
													30 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--14                             
													31 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--15 
													32 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--7
													33 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--8                  
													34 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--9	                                 
													35 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--10
													36 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--11
													37 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--12
													38 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--13
													39 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8)--14                              
													);
begin
--HANG 1
LCD_HANG_1(7 DOWNTO 0)			<= HOVATEN_TSP(0) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(0);
											
LCD_HANG_1(15 DOWNTO 8)			<= HOVATEN_TSP(1) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(1);
											
LCD_HANG_1(23 DOWNTO 16)		<= HOVATEN_TSP(2) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(2);
											
LCD_HANG_1(31 DOWNTO 24)		<= HOVATEN_TSP(3) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(3);

LCD_HANG_1(39 DOWNTO 32)		<= HOVATEN_TSP(4) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(4);

LCD_HANG_1(47 DOWNTO 40)		<= HOVATEN_TSP(5) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(5);

LCD_HANG_1(55 DOWNTO 48)		<= HOVATEN_TSP(6) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(6);

LCD_HANG_1(63 DOWNTO 56)		<= HOVATEN_TSP(7) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(7);

LCD_HANG_1(71 DOWNTO 64)		<= HOVATEN_TSP(8) WHEN CHOPHEP = '0' ELSE 
											HOVATEN_PST(8);

LCD_HANG_1(79 DOWNTO 72)		<= HOVATEN_TSP(9) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(9);

LCD_HANG_1(87 DOWNTO 80)		<= HOVATEN_TSP(10) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(10);

LCD_HANG_1(95 DOWNTO 88)		<= HOVATEN_TSP(11) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(11);

LCD_HANG_1(103 DOWNTO 96)		<= HOVATEN_TSP(12) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(12);

LCD_HANG_1(111 DOWNTO 104)		<= HOVATEN_TSP(13) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(13);

LCD_HANG_1(119 DOWNTO 112)		<= HOVATEN_TSP(14) WHEN CHOPHEP = '0' ELSE 
											HOVATEN_PST(14);
   	
LCD_HANG_1(127 DOWNTO 120)		<= HOVATEN_TSP(15) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(15);

LCD_HANG_1(135 DOWNTO 128) 	<= HOVATEN_TSP(16) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(16);

LCD_HANG_1(143 DOWNTO 136) 	<= HOVATEN_TSP(17) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(17);

LCD_HANG_1(151 DOWNTO 144) 	<= HOVATEN_TSP(18) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(18);

LCD_HANG_1(159 DOWNTO 152) 	<= HOVATEN_TSP(19) WHEN CHOPHEP = '0' ELSE
											HOVATEN_PST(19);



PROCESS(RST,ENA_DB,HOVATEN_TSP)
	 BEGIN
		IF (RST = '1') THEN 	HOVATEN_TSP <= (	0 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--19
															1 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('G'),8),--19
															2 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('Y'),8),--19
															3 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8),--19
															4 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--19
															5 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--19
															6 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('V'),8),--19
															7 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8),--16
															8 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--16
															9 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															10 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('V'),8),--16
															11 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('Y'),8),--16
															12 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															13 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															14 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															15 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															16 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															17 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--1
															18 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--2                              
															19 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--3                                   
															20 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--4
															21 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--5
															22 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--6
															23 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--7
															24 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--8                  
															25 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--9	                                 
															26 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--10
															27 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--11
															28 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--12
															29 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--13
															30 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--14                             
															31 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--15 
															32 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--7
															33 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--8                  
															34 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--9	                                 
															35 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--10
															36 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--11
															37 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--12
															38 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--13
															39 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8));
	ELSIF (FALLING_EDGE(ENA_DB)) THEN
		HOVATEN_TSP(39) <= HOVATEN_TSP(0);
		FOR I IN 0 TO 38
		LOOP
		 HOVATEN_TSP(I) <= HOVATEN_TSP(I+1);
		END LOOP;
	ELSE
		 HOVATEN_TSP <= HOVATEN_TSP;
	END IF;
END PROCESS;



PROCESS(RST,ENA_DB,HOVATEN_PST)
BEGIN
		IF (RST = '1') THEN 	HOVATEN_PST <= (	0 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--19
															1 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('G'),8),--19
															2 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('Y'),8),--19
															3 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8),--19
															4 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--19
															5 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--19
															6 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('V'),8),--19
															7 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8),--16
															8 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8),--16
															9 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															10 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('V'),8),--16
															11 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('Y'),8),--16
															12 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															13 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															14 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															15 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															16 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--16
															17 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--1
															18 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--2                              
															19 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--3                                   
															20 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--4
															21 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--5
															22 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--6
															23 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--7
															24 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--8                  
															25 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--9	                                 
															26 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--10
															27 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--11
															28 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--12
															29 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--13
															30 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--14                             
															31 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--15 
															32 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--7
															33 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--8                  
															34 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--9	                                 
															35 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--10
															36 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--11
															37 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--12
															38 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),--13
															39 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8));
	ELSIF (FALLING_EDGE(ENA_DB)) THEN
		HOVATEN_PST(0) <= HOVATEN_PST(39);
		FOR I IN 0 TO 38
		LOOP
		 HOVATEN_PST(I+1) <= HOVATEN_PST(I);
		END LOOP;
	ELSE
		 HOVATEN_PST <= HOVATEN_PST;
	END IF;
END PROCESS;

--HANG 2
LCD_HANG_2(7 DOWNTO 0) 			<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(15 DOWNTO 8) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(23 DOWNTO 16) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(31 DOWNTO 24) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(39 DOWNTO 32) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(47 DOWNTO 40) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(55 DOWNTO 48) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(63 DOWNTO 56) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(71 DOWNTO 64) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(79 DOWNTO 72) 		<= X"3" & CHUC;
LCD_HANG_2(87 DOWNTO 80) 		<= X"3" & DONVI;
LCD_HANG_2(95 DOWNTO 88) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(103 DOWNTO 96) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(111 DOWNTO 104) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(119 DOWNTO 112) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(127 DOWNTO 120) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(135 DOWNTO 128) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(143 DOWNTO 136) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(151 DOWNTO 144) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(159 DOWNTO 152) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);

---hang3
LCD_HANG_3(7 DOWNTO 0) 			<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(15 DOWNTO 8) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(23 DOWNTO 16) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(31 DOWNTO 24) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(39 DOWNTO 32) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(47 DOWNTO 40) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(55 DOWNTO 48) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(63 DOWNTO 56) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(71 DOWNTO 64) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(79 DOWNTO 72) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(87 DOWNTO 80) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(95 DOWNTO 88) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(103 DOWNTO 96) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(111 DOWNTO 104) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(119 DOWNTO 112) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(127 DOWNTO 120) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(135 DOWNTO 128) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(143 DOWNTO 136) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(151 DOWNTO 144) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_3(159 DOWNTO 152) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);

--hang4
LCD_HANG_4(7 DOWNTO 0) 			<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(15 DOWNTO 8) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(23 DOWNTO 16) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(31 DOWNTO 24) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(39 DOWNTO 32) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(47 DOWNTO 40) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(55 DOWNTO 48) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(63 DOWNTO 56) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(71 DOWNTO 64) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(79 DOWNTO 72) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(87 DOWNTO 80) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(95 DOWNTO 88) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(103 DOWNTO 96) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(111 DOWNTO 104) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(119 DOWNTO 112) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(127 DOWNTO 120) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(135 DOWNTO 128) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(143 DOWNTO 136) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(151 DOWNTO 144) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_4(159 DOWNTO 152) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);

end Behavioral;

