library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DEM_2SOB is
    Port ( CKHT,RST,ENA_DB,ENA_SS,ENA_SS1 : in  STD_LOGIC;
           DONVI,CHUC : out  STD_LOGIC_VECTOR (3 downto 0));
end DEM_2SOB;

architecture Behavioral of DEM_2SOB is
SIGNAL DONVI_REG, DONVI_NEXT: STD_LOGIC_VECTOR (3 DOWNTO 0):="0101";
SIGNAL CHUC_REG, CHUC_NEXT: STD_LOGIC_VECTOR (3 DOWNTO 0):= "0011";
begin
PROCESS (CKHT, RST)
	BEGIN
		IF RST ='1' OR CHUC_REG&DONVI_REG = "00100100" THEN DONVI_REG <= "0101";
							  CHUC_REG <= "0011";
		ELSIF FALLING_EDGE (CKHT) THEN DONVI_REG <= DONVI_NEXT;
													CHUC_REG <= CHUC_NEXT;
		END IF;
	END PROCESS;
--------------------------------------------------------------------
	PROCESS (DONVI_REG, CHUC_REG, ENA_SS, ENA_DB)
	BEGIN
		DONVI_NEXT <= DONVI_REG;
		CHUC_NEXT <= CHUC_REG;
		IF ENA_DB ='1' THEN 
			IF ENA_SS ='1' AND ENA_SS1 = '0' THEN 
					IF DONVI_REG /= X"0" THEN DONVI_NEXT <= DONVI_REG - 1;
					ELSE								
						DONVI_NEXT <= X"9";
						IF CHUC_REG /= X"0" THEN CHUC_NEXT <= CHUC_REG - 1;
						ELSE								
						CHUC_NEXT <= X"9";
						END IF;
					END IF;
			END IF;
		END IF;
	END PROCESS;
	DONVI <= DONVI_REG;
	CHUC <= CHUC_REG;
end Behavioral;



