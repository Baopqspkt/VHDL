
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE. STD_LOGIC_ARITH.ALL;


entity LCD_NHIET_DO_DS18B20 is
    Port ( CKHT: in  STD_LOGIC;
           BELL : out  STD_LOGIC;
			  BTN_N : in  STD_LOGIC_VECTOR (3 DOWNTO 0);
			  DS18B20 : inout  STD_LOGIC;
			  DECIMAL, LED : out  STD_LOGIC_VECTOR (3 downto 0);
           LCD_E, LCD_RS, LCD_RW : out  STD_LOGIC;
           LCD_DB : out  STD_LOGIC_VECTOR (7 downto 0));
end LCD_NHIET_DO_DS18B20;

architecture Behavioral of LCD_NHIET_DO_DS18B20 is

SIGNAL RST, DS_PRESENT,ENA5HZ,ENA10HZ,ENADB: STD_LOGIC;
SIGNAL DONVI, CHUC, TRAM,DVX,CHX: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL NHIETDO: STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL TEMPERATURE: STD_LOGIC_VECTOR (11 DOWNTO 0);
SIGNAL LCD_HANG_1: STD_LOGIC_VECTOR (159 DOWNTO 0);
SIGNAL LCD_HANG_2: STD_LOGIC_VECTOR (159 DOWNTO 0);
SIGNAL LCD_HANG_3: STD_LOGIC_VECTOR (159 DOWNTO 0);
SIGNAL LCD_HANG_4: STD_LOGIC_VECTOR (159 DOWNTO 0);
SIGNAL LED0, LED1, LED2: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL LCD_MA_DONVI:	STD_LOGIC_VECTOR (47 DOWNTO 0);
SIGNAL LCD_MA_CHUC:	STD_LOGIC_VECTOR (47 DOWNTO 0);
SIGNAL DV:	STD_LOGIC_VECTOR (47 DOWNTO 0);
SIGNAL CH:	STD_LOGIC_VECTOR (47 DOWNTO 0);
SIGNAL SEL1,SEL2,ENASS : STD_LOGIC;
begin

	LCD_RW <= '0';
	RST <= NOT BTN_N(0);
	
	NHIETDO <= TEMPERATURE (11 DOWNTO 4);
	DECIMAL <= TEMPERATURE (3 DOWNTO 0);

	
	BELL <= '1';
DS18B20_TEMPERATURE: ENTITY WORK.DS18B20_TEMPERATURE
	PORT MAP ( 	CKHT => CKHT,
					RST => RST,
					DS18B20 => DS18B20,
					DS_PRESENT => DS_PRESENT,
					TEMPERATURE_OUT => TEMPERATURE);
	PROCESS (DS_PRESENT, DONVI, CHUC, TRAM)
	BEGIN
		IF (DS_PRESENT = '0') THEN
									LED0 <= DONVI;
									LED1 <= CHUC;
									LED2 <= TRAM;
		ELSE
									LED0 <= X"E";
									LED1 <= X"E";
									LED2 <= X"E";
		END IF;
	END PROCESS;
	
	
HEXTOBCD: ENTITY WORK.HEXTOBCD_8BIT
			PORT MAP(	SOHEX8BIT => NHIETDO,
							DONVI => DONVI,
							CHUC => CHUC,
							TRAM => TRAM);	
-------------------------------------------------------							
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
			PORT MAP(	CKHT => CKHT,
							ENA5HZ => ENA5HZ,
							ENA10HZ => ENA10HZ);

--------------------------------------------------------
DEM_2SO:	ENTITY WORK.DEM_2SO
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_DB => ENA5HZ,
							ENA_SS => ENASS,
							DONVI => DVX,
							CHUC => CHX
							); -- THEM CHO NAY

									
LCD_GIAI_MA_SO_TO_DVX: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(SO_GIAI_MA => DVX,
				LCD_MA_TO => DV
					);
					
LCD_GIAI_MA_SO_TO_CHX: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP( 
				SO_GIAI_MA => CHX,
				LCD_MA_TO => CH
				);
DEM_1BIT_BTNSS: ENTITY WORK.DEM_1BIT_BTN
		PORT MAP(	CKHT => CKHT,
						RST => RST,
						BTN => NOT BTN_N(1),
						Q => ENASS);

DEM_1BIT_BTN1: ENTITY WORK.DEM_1BIT_BTN
		PORT MAP(	CKHT => CKHT,
						RST => RST,
						BTN => NOT BTN_N(2),
						Q => SEL1);
DEM_1BIT_BTN2: ENTITY WORK.DEM_1BIT_BTN
		PORT MAP(	CKHT => CKHT,
						RST => RST,
						BTN => NOT BTN_N(3),
						Q => SEL2);
						
LCD_GIAI_MA_SO_TO_DV: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(SO_GIAI_MA => LED0,
				LCD_MA_TO => LCD_MA_DONVI
					);
					
LCD_GIAI_MA_SO_TO_CH: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP( 
				SO_GIAI_MA => LED1,
				LCD_MA_TO => LCD_MA_CHUC
				);

					
LCD_GAN_DULIEU_1SO_TO: ENTITY WORK.LCD_GAN_DULIEU_1SO_TO
	PORT MAP(
				LCD_MA_DONVI => LCD_MA_DONVI,
				LCD_MA_CHUC => LCD_MA_CHUC,
				CH          => CH,
				DV          => DV,
				SEL1        => SEL1,
				SEL2        => SEL2,
				LCD_HANG_1 => LCD_HANG_1,
				LCD_HANG_2 => LCD_HANG_2,
				LCD_HANG_3 => LCD_HANG_3,
				LCD_HANG_4 => LCD_HANG_4);

LCD_KHOITAO_HIENTHI:	ENTITY WORK.LCD_KHOITAO_HIENTHI
		PORT MAP(	LCD_DB => LCD_DB,
						LCD_RS => LCD_RS,
						LCD_E => LCD_E,
						LCD_RST => RST,
						LCD_CK => CKHT,
						LCD_HANG_1 => LCD_HANG_1,
						LCD_HANG_2 => LCD_HANG_2,
						LCD_HANG_3 => LCD_HANG_3,
						LCD_HANG_4 => LCD_HANG_4);

end Behavioral;

