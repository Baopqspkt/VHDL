
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL; 


entity LCD_GAN_DULIEU_HIENTHI_3SO is
    Port ( 
				H1_13, H1_14, H1_15,H2_13, H2_14: IN STD_LOGIC_VECTOR (3 downto 0);
			  LCD_HANG_1 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_HANG_2 : out  STD_LOGIC_VECTOR (159 downto 0));
end LCD_GAN_DULIEU_HIENTHI_3SO;

architecture Behavioral of LCD_GAN_DULIEU_HIENTHI_3SO is
SIGNAL XOA: STD_LOGIC_VECTOR(3 DOWNTO 0);
begin
--HANG 1);
XOA <= H1_13;
LCD_HANG_1(7 DOWNTO 0) 			<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
LCD_HANG_1(15 DOWNTO 8) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
LCD_HANG_1(23 DOWNTO 16) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
LCD_HANG_1(31 DOWNTO 24) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
LCD_HANG_1(39 DOWNTO 32) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
LCD_HANG_1(47 DOWNTO 40) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_1(55 DOWNTO 48) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
LCD_HANG_1(63 DOWNTO 56) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
LCD_HANG_1(71 DOWNTO 64) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_1(79 DOWNTO 72) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
LCD_HANG_1(87 DOWNTO 80) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
LCD_HANG_1(95 DOWNTO 88) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
LCD_HANG_1(103 DOWNTO 96) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_1(111 DOWNTO 104) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_1(119 DOWNTO 112) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_1(127 DOWNTO 120) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8) WHEN XOA = "0000" ELSE X"3" & H1_13;
LCD_HANG_1(135 DOWNTO 128) 	<= X"3" & H1_14;
LCD_HANG_1(143 DOWNTO 136) 	<= X"3" & H1_15;
LCD_HANG_1(151 DOWNTO 144) 	<= X"00";
LCD_HANG_1(159 DOWNTO 152) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
--HANG 2
LCD_HANG_2(7 DOWNTO 0) 			<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
LCD_HANG_2(15 DOWNTO 8) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
LCD_HANG_2(23 DOWNTO 16) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
LCD_HANG_2(31 DOWNTO 24) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
LCD_HANG_2(39 DOWNTO 32) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
LCD_HANG_2(47 DOWNTO 40) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(55 DOWNTO 48) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
LCD_HANG_2(63 DOWNTO 56) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
LCD_HANG_2(71 DOWNTO 64) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(79 DOWNTO 72) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
LCD_HANG_2(87 DOWNTO 80) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
LCD_HANG_2(95 DOWNTO 88) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
LCD_HANG_2(103 DOWNTO 96) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
LCD_HANG_2(111 DOWNTO 104) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(119 DOWNTO 112) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(127 DOWNTO 120) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
LCD_HANG_2(135 DOWNTO 128) 	<= X"3" & H2_13;
LCD_HANG_2(143 DOWNTO 136) 	<= X"3" & H2_14;
LCD_HANG_2(151 DOWNTO 144) 	<= X"00";
LCD_HANG_2(159 DOWNTO 152) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
end Behavioral;

