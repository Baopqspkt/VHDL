library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity LCD_MR_HENTHI_DEM_LEN_XUONG_DICH_TSP_PST is
    Port ( CKHT : in  STD_LOGIC;
           BTN_N : in  STD_LOGIC_VECTOR (1 downto 0);
           BELL : out  STD_LOGIC;
           LCD_DB : out  STD_LOGIC_VECTOR (7 downto 0);
           LCD_RS : out  STD_LOGIC;
           LCD_RW : out  STD_LOGIC;
           LCD_E : out  STD_LOGIC);
end LCD_MR_HENTHI_DEM_LEN_XUONG_DICH_TSP_PST;

architecture Behavioral of LCD_MR_HENTHI_DEM_LEN_XUONG_DICH_TSP_PST is
SIGNAL RST:STD_LOGIC;
SIGNAL ENA_SS,ENA_DB:STD_LOGIC;
SIGNAL DONVI,CHUC:STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL LCD_HANG_1:STD_LOGIC_VECTOR(159 DOWNTO 0);
SIGNAL LCD_HANG_2:STD_LOGIC_VECTOR(159 DOWNTO 0);
SIGNAL LCD_HANG_3:STD_LOGIC_VECTOR(159 DOWNTO 0);
SIGNAL LCD_HANG_4:STD_LOGIC_VECTOR(159 DOWNTO 0);
SIGNAL CHOPHEP:STD_LOGIC;
begin

LCD_RW	<= '0';
BELL		<= '1';
RST		<= NOT BTN_N(0);


CHIA_10ENA:ENTITY WORK.CHIA_10ENA
PORT MAP (CKHT	=> CKHT,
			 ENA5HZ	=> ENA_DB);
			 
DEM_1BIT_BTN:ENTITY WORK.DEM_1BIT_BTN
PORT MAP( CKHT	=> CKHT,
			 BTN	=> NOT BTN_N(1),
			 RST	=> RST,
			 Q		=> ENA_SS);

DEM_2SO_UD:ENTITY WORK.DEM_2SO_UD
PORT MAP(ENA_DB	=> ENA_DB,
			CKHT		=> CKHT,
			RST		=> RST,
			ENA_SS	=> ENA_SS,
			ENA_UD	=> CHOPHEP,
			DONVI		=> DONVI,
			CHUC		=> CHUC);

LCD_GAN_DULIEU_HIENTHI_3_SO:ENTITY WORK.LCD_GAN_DULIEU_HIENTHI
PORT MAP ( DONVI	=> DONVI,
			  CHUC	=> CHUC,
			  RST		=> RST,
			  ENA_DB	=> ENA_DB,
			  CHOPHEP	=> CHOPHEP,
			  LCD_HANG_1	=> LCD_HANG_1,
			  LCD_HANG_2 	=> LCD_HANG_2,
			  LCD_HANG_3	=> LCD_HANG_3,
			  LCD_HANG_4 	=> LCD_HANG_4);

LCD_KHOITAO_HIENTHI:ENTITY WORK.LCD_KHOITAO_HIENTHI
PORT MAP (LCD_CK	=> CKHT,
			 LCD_RST	=> RST,
			 LCD_HANG_1	=> LCD_HANG_1,
			 LCD_HANG_2 => LCD_HANG_2,
			 LCD_HANG_3	=> LCD_HANG_3,
			 LCD_HANG_4 => LCD_HANG_4,
			 LCD_DB		=> LCD_DB,
			 LCD_E		=> LCD_E,
			 LCD_RS		=> LCD_RS);
			 
			 
end Behavioral;

