
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity LCD_DEM_00_99_SO_TO is
    Port ( CKHT, BTN_N0, SW0 : in  STD_LOGIC;
           BELL : out  STD_LOGIC;
           LCD_E, LCD_RS, LCD_RW : out  STD_LOGIC;
			  DS18B20 : inout  STD_LOGIC;
			  DECIMAL : out  STD_LOGIC_VECTOR (3 downto 0);
           LCD_DB : out  STD_LOGIC_VECTOR (7 downto 0)
			  );  
end LCD_DEM_00_99_SO_TO;

architecture Behavioral of LCD_DEM_00_99_SO_TO is
SIGNAL LCD_HANG_1	:	STD_LOGIC_VECTOR (159 downto 0);
SIGNAL LCD_HANG_2	:	STD_LOGIC_VECTOR (159 DOWNTO 0);
SIGNAL LCD_HANG_3	:	STD_LOGIC_VECTOR (159 downto 0);
SIGNAL LCD_HANG_4	:	STD_LOGIC_VECTOR (159 DOWNTO 0);

SIGNAL GIAY, PHUT, GIO: STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL GIO5: STD_LOGIC_VECTOR (4 DOWNTO 0);

SIGNAL CH_GIO, DV_GIO: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL CH_PHUT, DV_PHUT: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL CH_GIAY, DV_GIAY: STD_LOGIC_VECTOR (3 DOWNTO 0);

SIGNAL LCD_CH_GIO:	STD_LOGIC_VECTOR (47 DOWNTO 0);
SIGNAL LCD_DV_GIO:	STD_LOGIC_VECTOR (47 DOWNTO 0);

SIGNAL LCD_CH_PHUT:	STD_LOGIC_VECTOR (47 DOWNTO 0);
SIGNAL LCD_DV_PHUT:	STD_LOGIC_VECTOR (47 DOWNTO 0);

SIGNAL LCD_CH_GIAY:	STD_LOGIC_VECTOR (47 DOWNTO 0);
SIGNAL LCD_DV_GIAY:	STD_LOGIC_VECTOR (47 DOWNTO 0);

SIGNAL ENA,RST,ENA_DB,DS_PRESENT,OE : STD_LOGIC;
SIGNAL DV, CH,TR: STD_LOGIC_VECTOR (3 DOWNTO 0);

SIGNAL LCD_CH_ND:	STD_LOGIC_VECTOR (47 DOWNTO 0);
SIGNAL LCD_DV_ND:	STD_LOGIC_VECTOR (47 DOWNTO 0);
SIGNAL LCD_CHU_TO:	STD_LOGIC_VECTOR (47 DOWNTO 0);

SIGNAL DONVI, CHUC, TRAM: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL NHIETDO: STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL TEMPERATURE: STD_LOGIC_VECTOR (11 DOWNTO 0);

begin

	LCD_RW <= '0';
	RST <= NOT BTN_N0;
	BELL <= '1';

	NHIETDO <= TEMPERATURE (11 DOWNTO 4);
	DECIMAL <= TEMPERATURE (3 DOWNTO 0);
	
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
					PORT MAP( CKHT => CKHT,
								ENA5HZ => ENA_DB);
DEM_2SO:	ENTITY WORK.DEM_2SO
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_DB => ENA_DB,
							OE    => OE);
DEM_1BIT_BTN: ENTITY WORK.DEM_1BIT_BTN
		PORT MAP(	CKHT => CKHT,
						RST => RST,
						BTN => OE,
						Q => ENA);

DS18B20_TEMPERATURE: ENTITY WORK.DS18B20_TEMPERATURE
	PORT MAP ( 	CKHT => CKHT,
					RST => RST,
					DS18B20 => DS18B20,
					DS_PRESENT => DS_PRESENT,
					TEMPERATURE_OUT => TEMPERATURE);
					
	PROCESS (DS_PRESENT, DONVI, CHUC, TRAM)
	BEGIN
		IF (DS_PRESENT = '0') THEN
									DV <= DONVI;
									CH <= CHUC;
									TR <= TRAM;
		ELSE
									DV <= X"E";
									CH <= X"E";
									TR <= X"E";
		END IF;
	END PROCESS;
	
	
HEXTOBCD: ENTITY WORK.HEXTOBCD_8BIT
			PORT MAP(	SOHEX8BIT => NHIETDO,
							DONVI => DONVI,
							CHUC => CHUC,
							TRAM => TRAM);		
----------------------------------------------------------------------------------------						
LCD_GIAI_MA_SO_TO_DV: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP( 
				SO_GIAI_MA => DV,
				LCD_MA_TO => LCD_DV_ND
				);
					
LCD_GIAI_MA_SO_TO_CH: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP( 
				SO_GIAI_MA => CH,
				LCD_MA_TO => LCD_CH_ND
				); 
								
DEM_GIOPHUTGIAY: ENTITY WORK.DEM_GIOPHUTGIAY
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_DB => ENA_DB,
							GIO => GIO5,
							PHUT => PHUT,
							GIAY => GIAY);
							
HEXTOBCD_GIO: ENTITY WORK.HEXTOBCD_6BIT
			PORT MAP(	SOHEX6BIT => GIO,
							DONVI => DV_GIO,
							CHUC => CH_GIO);
							
HEXTOBCD_PHUT: ENTITY WORK.HEXTOBCD_6BIT
			PORT MAP(	SOHEX6BIT => PHUT,
							DONVI => DV_PHUT,
							CHUC => CH_PHUT);
							
HEXTOBCD_GIAY: ENTITY WORK.HEXTOBCD_6BIT
			PORT MAP(	SOHEX6BIT => GIAY,
							DONVI => DV_GIAY,
							CHUC => CH_GIAY);	
LCD_GIAI_MA_SO_TO_CH_GIO: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(SO_GIAI_MA => CH_GIO,
				LCD_MA_TO => LCD_CH_GIO);
					
LCD_GIAI_MA_SO_TO_DV_GIO: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(SO_GIAI_MA => DV_GIO,
				LCD_MA_TO => LCD_DV_GIO);		
			
LCD_GIAI_MA_SO_TO_CH_PHUT: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(SO_GIAI_MA => CH_PHUT,
				LCD_MA_TO => LCD_CH_PHUT);
					
LCD_GIAI_MA_SO_TO_DV_PHUT: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(SO_GIAI_MA => DV_PHUT,
				LCD_MA_TO => LCD_DV_PHUT);		

LCD_GIAI_MA_CHU_TO: ENTITY WORK.LCD_GIAI_MA_CHU_TO
	PORT MAP(SO_GIAI_MA => X"C",
				LCD_MA_TO => LCD_CHU_TO);	

LCD_GIAI_MA_SO_TO_CH_GIAY: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(SO_GIAI_MA => CH_GIAY,
				LCD_MA_TO => LCD_CH_GIAY);
					
LCD_GIAI_MA_SO_TO_DV_GIAY: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(SO_GIAI_MA => DV_GIAY,
				LCD_MA_TO => LCD_DV_GIAY);					
LCD_GAN_DULIEU_1SO_TO: ENTITY WORK.LCD_GAN_DULIEU_1SO_TO
PORT MAP(
				CH_GIO	=> CH_GIO,
				DV_GIO	=> DV_GIO,
				
				CH_ND	=> CH,
				DV_ND	=> DV,
				
				CH_PHUT => CH_PHUT,
				DV_PHUT	=> DV_PHUT,
				
				CH_GIAY	=> CH_GIAY,
				DV_GIAY => DV_GIAY,
				
				LCD_CH_GIO => LCD_CH_GIO,
				LCD_DV_GIO => LCD_DV_GIO,
				LCD_CH_PHUT => LCD_CH_PHUT,
				LCD_DV_PHUT => LCD_DV_PHUT,
				LCD_CH_GIAY => LCD_CH_GIAY,
				LCD_DV_GIAY => LCD_DV_GIAY,
				LCD_CH_ND => LCD_CH_ND,
				LCD_DV_ND => LCD_DV_ND,
				LCD_CHU_TO => LCD_CHU_TO,
				
				ENA        => ENA,
				LCD_HANG_1 => LCD_HANG_1,
				LCD_HANG_2 => LCD_HANG_2,
				LCD_HANG_3 => LCD_HANG_3,
				LCD_HANG_4 => LCD_HANG_4);

LCD_KHOITAO_HIENTHI_CGRAM_SO_TO: ENTITY WORK.LCD_KHOITAO_HIENTHI_CGRAM_SO_TO
	PORT MAP(
				LCD_DB => LCD_DB,
				LCD_RS => LCD_RS,
				LCD_E => LCD_E,
				LCD_RST => RST,
				LCD_CK => CKHT,
				ENA    => ENA,
				LCD_HANG_1 => LCD_HANG_1,
				LCD_HANG_2 => LCD_HANG_2,
				LCD_HANG_3 => LCD_HANG_3,
				LCD_HANG_4 => LCD_HANG_4);
end Behavioral;

